package definitions;

parameter OPCODE_BRANCH = 7'h63;
parameter OPCODE_JALR   = 7'h67;
parameter OPCODE_JAL    = 7'h6f;
parameter OPCODE_OPIMM  = 7'h13;
parameter OPCODE_OP     = 7'h33;
parameter OPCODE_LOAD   = 7'h03;
parameter OPCODE_STORE  = 7'h23;

parameter ALU_
